-- ROM-based tile memory
library ieee;
